module TLcontroller(
    
    );
endmodule